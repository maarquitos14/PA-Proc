module cache(input clk, input rst, input [31:0] addr, output [31:0] data);
	assign data = 32'hffffffff;
endmodule 